module andgate (
input logic a,
input logic b,
output logic f
);
and u_and(f, a, b); // AND gate
endmodule
